`timescale 1ns/1ns

module ALU_Control (

);

endmodule