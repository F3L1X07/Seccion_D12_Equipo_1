`timescale 1ns/1ns

module Unidad_Control (
    //Entradas
    input [31:26]Instruccion,

    //Salidas
    output RegDst,
    output Branch,
    output MemRead,
    output MemtoReg,
    output ALUOp,
    output MemWrite,
    output ALUSrc,
    output RegWrite
);



endmodule