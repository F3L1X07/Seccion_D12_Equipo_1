`timescale 1ns/1ns

module MUX (

);

endmodule
