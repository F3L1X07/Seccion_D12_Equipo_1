`timescale 1ns/1ns

module Add_1 (
    //Entradas
    input PC_In,
    input CONST,

    //Salidas
    output Res
);

CONST = 4'd4;

endmodule
