`timescale 1ns/1ns

module Instruct_Memory (

);

endmodule
