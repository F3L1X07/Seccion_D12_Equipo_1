`timescale 1ns/1ns

module PC (
    //Entradas
    input [31:0]A,
    input CLK,

    //Salidas
    output [31:0]S
);

always @(posedge clk)     
begin                                                     
    salida = entrada
end

endmodule
