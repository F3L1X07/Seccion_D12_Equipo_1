`timescale 1ns/1ns

module Unidad_Control (

);

endmodule