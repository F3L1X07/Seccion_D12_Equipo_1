`timescale 1ns/1ns

module Instruction_Memory (

);

endmodule
