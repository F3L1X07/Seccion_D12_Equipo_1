`timescale 1ns/1ns

module Add_1 (
    //Entradas
    input PC_In,
    input [3:0]CONST,

    //Salidas
    output Res
);

assign CONST = 4'd4;

endmodule
