`timescale 1ns/1ns

module Banco_Registro (
    //Inputs
    input 
    
    //Outputs
    output 
);

endmodule